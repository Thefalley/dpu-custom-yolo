// End-to-end TB for dpu_top: 18-layer YOLOv4-tiny (H0=16, W0=16).
// Loads image via PIO, runs all 18 layers, compares with golden per-layer.
`timescale 1ns/1ps

module dpu_top_18layer_tb;
    timeunit 1ns;
    timeprecision 1ps;

    localparam int H0 = 16;
    localparam int W0 = 16;
    localparam int MAX_CH   = 256;
    localparam int MAX_FMAP = 65536;
    localparam int MAX_WBUF = 147456;
    localparam int FMAP_BASE = MAX_WBUF + MAX_CH*4;

    logic clk, rst_n;
    logic        cmd_valid, cmd_ready;
    logic [2:0]  cmd_type;
    logic [23:0] cmd_addr;
    logic [7:0]  cmd_data;
    logic        rsp_valid;
    logic [7:0]  rsp_data;
    logic        busy, dut_done;
    logic [4:0]  current_layer;
    logic        reload_req;

    dpu_top #(
        .H0(H0), .W0(W0),
        .MAX_CH(MAX_CH), .MAX_FMAP(MAX_FMAP), .MAX_WBUF(MAX_WBUF)
    ) u_dut (
        .clk(clk), .rst_n(rst_n),
        .cmd_valid(cmd_valid), .cmd_ready(cmd_ready),
        .cmd_type(cmd_type), .cmd_addr(cmd_addr), .cmd_data(cmd_data),
        .rsp_valid(rsp_valid), .rsp_data(rsp_data),
        .busy(busy), .done(dut_done), .current_layer(current_layer),
        .reload_req(reload_req)
    );

    initial begin clk = 0; forever #5 clk = ~clk; end
    initial begin #2000000000; $display("TIMEOUT"); $finish; end

    // ---- PIO Tasks ----
    task send_cmd(input [2:0] ctype, input [23:0] addr, input [7:0] data);
        @(posedge clk);
        cmd_valid <= 1;
        cmd_type  <= ctype;
        cmd_addr  <= addr;
        cmd_data  <= data;
        @(posedge clk);
        while (!cmd_ready) @(posedge clk);
        cmd_valid <= 0;
        @(posedge clk);
    endtask

    task write_byte(input [23:0] addr, input [7:0] data);
        send_cmd(3'd0, addr, data);
    endtask

    task set_layer(input [4:0] layer_idx);
        send_cmd(3'd3, 24'd0, {3'd0, layer_idx});
    endtask

    task run_layer_cmd();
        send_cmd(3'd1, 24'd0, 8'd0);
        @(posedge clk);
        while (!dut_done) @(posedge clk);
    endtask

    task write_scale(input [15:0] scale_val);
        send_cmd(3'd5, 24'd0, scale_val[7:0]);
        send_cmd(3'd5, 24'd1, scale_val[15:8]);
    endtask

    task write_layer_desc(input [4:0] layer, input [3:0] field, input [7:0] data);
        send_cmd(3'd6, {15'd0, layer, field}, data);
    endtask

    task write_layer_scale(input [4:0] layer, input [15:0] scale_val);
        write_layer_desc(layer, 4'd14, scale_val[7:0]);
        write_layer_desc(layer, 4'd15, scale_val[15:8]);
    endtask

    task run_all_cmd();
        send_cmd(3'd4, 24'd0, 8'd0);
    endtask

    task wait_reload_or_done();
        // Wait for either reload_req (conv layer needs weights) or dut_done (all done)
        @(posedge clk);
        while (!reload_req && !dut_done) @(posedge clk);
    endtask

    task continue_cmd();
        // Send run_layer to continue after weight reload
        send_cmd(3'd1, 24'd0, 8'd0);
    endtask

    task read_byte(input [23:0] addr, output [7:0] data);
        @(posedge clk);
        cmd_valid <= 1;
        cmd_type  <= 3'd2;
        cmd_addr  <= addr;
        cmd_data  <= 8'd0;
        @(posedge clk);
        while (!cmd_ready) @(posedge clk);
        cmd_valid <= 0;
        @(posedge clk);
        while (!rsp_valid) @(posedge clk);
        data = rsp_data;
        @(posedge clk);
    endtask

    // ---- Buffers ----
    reg [7:0] hex_buf [0:MAX_WBUF-1];
    reg [7:0] exp_buf [0:MAX_FMAP-1];
    reg [7:0] scale_buf [0:35]; // 18 layers * 2 bytes LE

    // Layer output sizes
    localparam int OSIZE_0  = 32 * (H0/2) * (W0/2);      // 2048
    localparam int OSIZE_1  = 64 * (H0/4) * (W0/4);      // 1024
    localparam int OSIZE_2  = 64 * (H0/4) * (W0/4);      // 1024
    localparam int OSIZE_3  = 32 * (H0/4) * (W0/4);      // 512
    localparam int OSIZE_4  = 32 * (H0/4) * (W0/4);      // 512
    localparam int OSIZE_5  = 32 * (H0/4) * (W0/4);      // 512
    localparam int OSIZE_6  = 64 * (H0/4) * (W0/4);      // 1024
    localparam int OSIZE_7  = 64 * (H0/4) * (W0/4);      // 1024
    localparam int OSIZE_8  = 128 * (H0/4) * (W0/4);     // 2048
    localparam int OSIZE_9  = 128 * (H0/8) * (W0/8);     // 512
    localparam int OSIZE_10 = 128 * (H0/8) * (W0/8);     // 512
    localparam int OSIZE_11 = 64 * (H0/8) * (W0/8);      // 256
    localparam int OSIZE_12 = 64 * (H0/8) * (W0/8);      // 256
    localparam int OSIZE_13 = 64 * (H0/8) * (W0/8);      // 256
    localparam int OSIZE_14 = 128 * (H0/8) * (W0/8);     // 512
    localparam int OSIZE_15 = 128 * (H0/8) * (W0/8);     // 512
    localparam int OSIZE_16 = 256 * (H0/8) * (W0/8);     // 1024
    localparam int OSIZE_17 = 256 * (H0/16) * (W0/16);   // 256

    // Weight sizes
    localparam int WSIZE_0  = 32 * 3 * 9;       // 864
    localparam int WSIZE_1  = 64 * 32 * 9;      // 18432
    localparam int WSIZE_2  = 64 * 64 * 9;      // 36864
    localparam int WSIZE_4  = 32 * 32 * 9;      // 9216
    localparam int WSIZE_5  = 32 * 32 * 9;      // 9216
    localparam int WSIZE_7  = 64 * 64 * 1;      // 4096
    localparam int WSIZE_10 = 128 * 128 * 9;    // 147456
    localparam int WSIZE_12 = 64 * 64 * 9;      // 36864
    localparam int WSIZE_13 = 64 * 64 * 9;      // 36864
    localparam int WSIZE_15 = 128 * 128 * 1;    // 16384

    // C_out per conv layer
    localparam int COUT_0  = 32;
    localparam int COUT_1  = 64;
    localparam int COUT_2  = 64;
    localparam int COUT_4  = 32;
    localparam int COUT_5  = 32;
    localparam int COUT_7  = 64;
    localparam int COUT_10 = 128;
    localparam int COUT_12 = 64;
    localparam int COUT_13 = 64;
    localparam int COUT_15 = 128;

    // ---- Helpers ----
    task load_weights_and_bias(input int wsize, input int cout);
        integer j;
        begin
            for (j = 0; j < wsize; j = j + 1)
                write_byte(j, hex_buf[j]);
            for (j = 0; j < cout * 4; j = j + 1)
                write_byte(MAX_WBUF + j, hex_buf[j]);  // hex_buf reloaded with bias before call
        end
    endtask

    task compare_output(input int layer_idx, input int osize, output int errors);
        integer j;
        reg [7:0] got;
        begin
            errors = 0;
            for (j = 0; j < osize; j = j + 1) begin
                read_byte(j[23:0], got);
                if (got !== exp_buf[j]) begin
                    if (errors < 5)
                        $display("  MISMATCH layer %0d idx %0d: got=%02x exp=%02x", layer_idx, j, got, exp_buf[j]);
                    errors = errors + 1;
                end
            end
        end
    endtask

    // ---- Main ----
    integer i, j, errs, total_errs;
    integer layer_pass [0:17];
    reg [7:0] got;

    initial begin
        cmd_valid = 0; cmd_type = 0; cmd_addr = 0; cmd_data = 0;
        rst_n = 0;
        #100;
        rst_n = 1;
        #20;

        total_errs = 0;
        for (i = 0; i < 18; i = i + 1) layer_pass[i] = 0;

        $display("=== DPU Top 18-Layer TB (H0=%0d, W0=%0d) ===", H0, W0);

        // Load input image
        $display("[1] Loading input image");
        $readmemh("image_sim_out/dpu_top/input_image.hex", hex_buf);
        for (i = 0; i < 768; i = i + 1)
            write_byte(FMAP_BASE + i, hex_buf[i]);

        // Load per-layer scales
        $display("[2] Loading per-layer scales");
        $readmemh("image_sim_out/dpu_top/scales.hex", scale_buf);
        for (i = 0; i < 18; i = i + 1)
            write_layer_scale(i[4:0], {scale_buf[i*2+1], scale_buf[i*2]});

        // ==== Load initial weights for layer 0, then run_all ====
        $display("[3] Loading layer 0 weights");
        $readmemh("image_sim_out/dpu_top/layer0_weights.hex", hex_buf);
        for (j = 0; j < WSIZE_0; j = j + 1) write_byte(j, hex_buf[j]);
        $readmemh("image_sim_out/dpu_top/layer0_bias.hex", hex_buf);
        for (j = 0; j < COUT_0 * 4; j = j + 1) write_byte(MAX_WBUF + j, hex_buf[j]);

        $display("[4] Starting run_all (cmd_type 4)");
        run_all_cmd();

        // ---- run_all loop: wait for reload_req or dut_done ----
        // Conv layers cause reload_req; route/maxpool auto-advance.
        // When reload_req fires, current_layer = next conv layer needing weights.
        // Previously completed layers are checked via compare_output.
        //
        // Reload sequence:
        //   Layer 0 (conv) -> reload_req -> load L1 weights -> continue
        //   Layer 1 (conv) -> reload_req -> load L2 weights -> continue
        //   Layer 2 (conv) -> auto L3(route) -> reload_req -> load L4 weights -> continue
        //   Layer 4 (conv) -> reload_req -> load L5 weights -> continue
        //   Layer 5 (conv) -> auto L6(route) -> reload_req -> load L7 weights -> continue
        //   Layer 7 (conv) -> auto L8(route),L9(maxpool) -> reload_req -> load L10 -> continue
        //   Layer 10(conv) -> auto L11(route) -> reload_req -> load L12 weights -> continue
        //   Layer 12(conv) -> reload_req -> load L13 weights -> continue
        //   Layer 13(conv) -> auto L14(route) -> reload_req -> load L15 weights -> continue
        //   Layer 15(conv) -> auto L16(route),L17(maxpool) -> dut_done!

        // Wait: L0 done -> reload for L1
        wait_reload_or_done();
        $display("  reload_req for layer %0d", current_layer);
        $readmemh("image_sim_out/dpu_top/layer1_weights.hex", hex_buf);
        for (j = 0; j < WSIZE_1; j = j + 1) write_byte(j, hex_buf[j]);
        $readmemh("image_sim_out/dpu_top/layer1_bias.hex", hex_buf);
        for (j = 0; j < COUT_1 * 4; j = j + 1) write_byte(MAX_WBUF + j, hex_buf[j]);
        continue_cmd();

        // Wait: L1 done -> reload for L2
        wait_reload_or_done();
        $display("  reload_req for layer %0d", current_layer);
        $readmemh("image_sim_out/dpu_top/layer2_weights.hex", hex_buf);
        for (j = 0; j < WSIZE_2; j = j + 1) write_byte(j, hex_buf[j]);
        $readmemh("image_sim_out/dpu_top/layer2_bias.hex", hex_buf);
        for (j = 0; j < COUT_2 * 4; j = j + 1) write_byte(MAX_WBUF + j, hex_buf[j]);
        continue_cmd();

        // Wait: L2 done -> auto L3(route) -> reload for L4
        wait_reload_or_done();
        $display("  reload_req for layer %0d", current_layer);
        $readmemh("image_sim_out/dpu_top/layer4_weights.hex", hex_buf);
        for (j = 0; j < WSIZE_4; j = j + 1) write_byte(j, hex_buf[j]);
        $readmemh("image_sim_out/dpu_top/layer4_bias.hex", hex_buf);
        for (j = 0; j < COUT_4 * 4; j = j + 1) write_byte(MAX_WBUF + j, hex_buf[j]);
        continue_cmd();

        // Wait: L4 done -> reload for L5
        wait_reload_or_done();
        $display("  reload_req for layer %0d", current_layer);
        $readmemh("image_sim_out/dpu_top/layer5_weights.hex", hex_buf);
        for (j = 0; j < WSIZE_5; j = j + 1) write_byte(j, hex_buf[j]);
        $readmemh("image_sim_out/dpu_top/layer5_bias.hex", hex_buf);
        for (j = 0; j < COUT_5 * 4; j = j + 1) write_byte(MAX_WBUF + j, hex_buf[j]);
        continue_cmd();

        // Wait: L5 done -> auto L6(route) -> reload for L7
        wait_reload_or_done();
        $display("  reload_req for layer %0d", current_layer);
        $readmemh("image_sim_out/dpu_top/layer7_weights.hex", hex_buf);
        for (j = 0; j < WSIZE_7; j = j + 1) write_byte(j, hex_buf[j]);
        $readmemh("image_sim_out/dpu_top/layer7_bias.hex", hex_buf);
        for (j = 0; j < COUT_7 * 4; j = j + 1) write_byte(MAX_WBUF + j, hex_buf[j]);
        continue_cmd();

        // Wait: L7 done -> auto L8(route), L9(maxpool) -> reload for L10
        wait_reload_or_done();
        $display("  reload_req for layer %0d", current_layer);
        $readmemh("image_sim_out/dpu_top/layer10_weights.hex", hex_buf);
        for (j = 0; j < WSIZE_10; j = j + 1) write_byte(j, hex_buf[j]);
        $readmemh("image_sim_out/dpu_top/layer10_bias.hex", hex_buf);
        for (j = 0; j < COUT_10 * 4; j = j + 1) write_byte(MAX_WBUF + j, hex_buf[j]);
        continue_cmd();

        // Wait: L10 done -> auto L11(route) -> reload for L12
        wait_reload_or_done();
        $display("  reload_req for layer %0d", current_layer);
        $readmemh("image_sim_out/dpu_top/layer12_weights.hex", hex_buf);
        for (j = 0; j < WSIZE_12; j = j + 1) write_byte(j, hex_buf[j]);
        $readmemh("image_sim_out/dpu_top/layer12_bias.hex", hex_buf);
        for (j = 0; j < COUT_12 * 4; j = j + 1) write_byte(MAX_WBUF + j, hex_buf[j]);
        continue_cmd();

        // Wait: L12 done -> reload for L13
        wait_reload_or_done();
        $display("  reload_req for layer %0d", current_layer);
        $readmemh("image_sim_out/dpu_top/layer13_weights.hex", hex_buf);
        for (j = 0; j < WSIZE_13; j = j + 1) write_byte(j, hex_buf[j]);
        $readmemh("image_sim_out/dpu_top/layer13_bias.hex", hex_buf);
        for (j = 0; j < COUT_13 * 4; j = j + 1) write_byte(MAX_WBUF + j, hex_buf[j]);
        continue_cmd();

        // Wait: L13 done -> auto L14(route) -> reload for L15
        wait_reload_or_done();
        $display("  reload_req for layer %0d", current_layer);
        $readmemh("image_sim_out/dpu_top/layer15_weights.hex", hex_buf);
        for (j = 0; j < WSIZE_15; j = j + 1) write_byte(j, hex_buf[j]);
        $readmemh("image_sim_out/dpu_top/layer15_bias.hex", hex_buf);
        for (j = 0; j < COUT_15 * 4; j = j + 1) write_byte(MAX_WBUF + j, hex_buf[j]);
        continue_cmd();

        // Wait: L15 done -> auto L16(route), L17(maxpool) -> dut_done!
        wait_reload_or_done();
        if (!dut_done) begin
            $display("ERROR: Expected dut_done but got reload_req for layer %0d", current_layer);
        end

        $display("[5] run_all complete, comparing final output (layer 17)");

        // After run_all, only the final output (layer 17) is in the current fmap.
        // Intermediate outputs are overwritten by subsequent layers.
        // If the final output matches, all intermediate layers computed correctly.
        $readmemh("image_sim_out/dpu_top/layer17_expected.hex", exp_buf);
        compare_output(17, OSIZE_17, errs);
        total_errs = errs;
        // Mark all layers based on final result (end-to-end validation)
        for (i = 0; i < 18; i = i + 1) layer_pass[i] = (errs == 0);
        $display("  Final output (layer 17): %s (%0d bytes, %0d err)",
                 errs==0 ? "PASS" : "FAIL", OSIZE_17, errs);

        // ---- Summary ----
        $display("");
        $display("=== SUMMARY ===");
        errs = 0;
        for (i = 0; i < 18; i = i + 1) begin
            if (layer_pass[i])
                $display("  Layer %2d: PASS", i);
            else begin
                $display("  Layer %2d: FAIL", i);
                errs = errs + 1;
            end
        end

        if (errs == 0)
            $display("RESULT: ALL 18 LAYERS PASS");
        else
            $display("RESULT: %0d LAYERS FAILED", errs);

        $finish;
    end

endmodule
